module adder (Reset, clk, A, B, computerPress);

	input logic Reset, clk;
	
	input logic [9:0] A, B;
	
	output logic computerPress;
	
	
